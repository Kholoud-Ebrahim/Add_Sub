package add_sub_pkg;
    import uvm_pkg::*;
    import param_pkg::*;
    `include "uvm_macros.svh"
     
    `include "add_sequence_item.svh"
    `include "sub_sequence_item.svh"

    `include "add_base_sequence.svh"    
    `include "sub_base_sequence.svh"    
    `include "add_full_sequence.svh"    
    `include "sub_full_sequence.svh"    
    `include "add_null_sequence.svh"    
    `include "sub_null_sequence.svh"    
  
    `include "add_sequencer.svh"
    `include "sub_sequencer.svh"

    `include "add_driver.svh"   
    `include "sub_driver.svh"

    `include "add_monitor.svh"   
    `include "sub_monitor.svh"   

    `include "add_agent.svh"  
    `include "sub_agent.svh"   

    `include "add_scoreboard.svh"  
    `include "sub_scoreboard.svh"   
    
    `include "add_sub_env.svh"  

    `include "add_sub_base_test.svh"
    `include "add_sub_fulls_test.svh" 
    `include "add_sub_nulls_test.svh" 
    `include "add_sub_random_test.svh" 

endpackage :add_sub_pkg