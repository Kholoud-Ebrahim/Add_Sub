package param_pkg;
    parameter WIDTH = 10;
    parameter CLK_PERIOD = 20ns;
endpackage :param_pkg